-- 31 x 31 px

constant ZERO: char:= (
				"0000000000000000000000000000000",
				"0000000000000111110000000000000",
				"0000000000001111111000000000000",
				"0000000000011110111100000000000",
				"0000000000111100011110000000000",
				"0000000001111100011111000000000",
				"0000000001111100011111000000000",
				"0000000001111100011111000000000",
				"0000000011111100011111100000000",
				"0000000011111100011111100000000",
				"0000000011111100011111100000000",
				"0000000011111100011111100000000",
				"0000000011111100011111100000000",
				"0000000011111100011111100000000",
				"0000000111111100011111110000000",
				"0000000111111100011111110000000",
				"0000000111111100011111110000000",
				"0000000011111100011111100000000",
				"0000000011111100011111100000000",
				"0000000011111100011111100000000",
				"0000000011111100011111100000000",
				"0000000011111100011111100000000",
				"0000000011111100011111100000000",
				"0000000011111100011111100000000",
				"0000000001111100011111000000000",
				"0000000001111100011111000000000",
				"0000000000111100011110000000000",
				"0000000000111100011110000000000",
				"0000000000011111111100000000000",
				"0000000000001111110000000000000",
				"0000000000000000000000000000000"
					);
					
constant ONE: char:= (
				"0000000000000000000000000000000",
				"0000000000000000011000000000000",
				"0000000000000000111000000000000",
				"0000000000000001111000000000000",
				"0000000000000011111000000000000",
				"0000000000000111111000000000000",
				"0000000000001111111000000000000",
				"0000000000111111111000000000000",
				"0000000000111111111000000000000",
				"0000000000000111111000000000000",
				"0000000000000111111000000000000",
				"0000000000000111111000000000000",
				"0000000000000111111000000000000",
				"0000000000000111111000000000000",
				"0000000000000111111000000000000",
				"0000000000000111111000000000000",
				"0000000000000111111000000000000",
				"0000000000000111111000000000000",
				"0000000000000111111000000000000",
				"0000000000000111111000000000000",
				"0000000000000111111000000000000",
				"0000000000000111111000000000000",
				"0000000000000111111000000000000",
				"0000000000000111111000000000000",
				"0000000000000111111000000000000",
				"0000000000000111111000000000000",
				"0000000000000111111000000000000",
				"0000000000000111111100000000000",
				"0000000000011111111110000000000",
				"0000000000011111111110000000000",
				"0000000000000000000000000000000"
					);

constant TWO: char:= (
				"0000000000000000000000000000000",
				"0000000000001111110000000000000",
				"0000000000111111111100000000000",
				"0000000001111101111110000000000",
				"0000000001111000111111000000000",
				"0000000011111000011111100000000",
				"0000000011111000011111100000000",
				"0000000011111000011111100000000",
				"0000000011111000011111100000000",
				"0000000011111000011111100000000",
				"0000000001110000011111100000000",
				"0000000000000000011111100000000",
				"0000000000000000111111100000000",
				"0000000000000000111111000000000",
				"0000000000000000111111000000000",
				"0000000000000001111110000000000",
				"0000000000000001111100000000000",
				"0000000000000011111000000000000",
				"0000000000000111110000000000000",
				"0000000000001111100000000000000",
				"0000000000001110000000000000000",
				"0000000000011100000000000000000",
				"0000000000111000000001110000000",
				"0000000001110000000001100000000",
				"0000000011100000000001100000000",
				"0000000011111111111111100000000",
				"0000000011111111111111100000000",
				"0000000111111111111111100000000",
				"0000000111111111111111100000000",
				"0000000111111111111111000000000",
				"0000000000000000000000000000000"
					);

constant THREE: char:= (
				"0000000000000000000000000000000",
				"0000000000011111110000000000000",
				"0000000001111111111000000000000",
				"0000000001110001111100000000000",
				"0000000011110001111110000000000",
				"0000000011110001111110000000000",
				"0000000111110001111111000000000",
				"0000000111110001111111000000000",
				"0000000011110001111111000000000",
				"0000000011110001111111000000000",
				"0000000000000001111110000000000",
				"0000000000000001111110000000000",
				"0000000000000001111100000000000",
				"0000000000011111111000000000000",
				"0000000000111111100000000000000",
				"0000000000111111111000000000000",
				"0000000000000001111100000000000",
				"0000000000000001111110000000000",
				"0000000000000000111111000000000",
				"0000000000000000111111000000000",
				"0000000000000000111111000000000",
				"0000000011100000111111100000000",
				"0000000111110000111111100000000",
				"0000000111110000111111100000000",
				"0000000111110000111111000000000",
				"0000000111110000111111000000000",
				"0000000011110000111110000000000",
				"0000000011110001111110000000000",
				"0000000001111111111100000000000",
				"0000000000111111110000000000000",
				"0000000000000000000000000000000"
					);

constant FOUR: char:= (
				"0000000000000000000000000000000",
				"0000000000000000011100000000000",
				"0000000000000000011100000000000",
				"0000000000000000111100000000000",
				"0000000000000000111100000000000",
				"0000000000000001111100000000000",
				"0000000000000011111100000000000",
				"0000000000000011111100000000000",
				"0000000000000111111100000000000",
				"0000000000001111111100000000000",
				"0000000000001111111100000000000",
				"0000000000011111111100000000000",
				"0000000000011011111100000000000",
				"0000000000111011111100000000000",
				"0000000001110011111100000000000",
				"0000000001100011111100000000000",
				"0000000011100011111100000000000",
				"0000000011000011111100000000000",
				"0000000110000011111100000000000",
				"0000001110000011111100000000000",
				"0000001111111111111111100000000",
				"0000001111111111111111100000000",
				"0000000111111111111111000000000",
				"0000000000000011111100000000000",
				"0000000000000011111100000000000",
				"0000000000000011111100000000000",
				"0000000000000011111100000000000",
				"0000000000000011111110000000000",
				"0000000000000111111111000000000",
				"0000000000000111111111000000000",
				"0000000000000000000000000000000"
					);

constant FIVE: char:= (
				"0000000000000000000110000000000",
				"0000000000111111111110000000000",
				"0000000000111111111110000000000",
				"0000000000111111111110000000000",
				"0000000000111111111110000000000",
				"0000000000111111111110000000000",
				"0000000000110000000000000000000",
				"0000000001110000000000000000000",
				"0000000001110000000000000000000",
				"0000000001100000000000000000000",
				"0000000001100001000000000000000",
				"0000000001111111111000000000000",
				"0000000001111111111100000000000",
				"0000000001110001111110000000000",
				"0000000001110000111111000000000",
				"0000000001100000111111000000000",
				"0000000000000000111111100000000",
				"0000000000000000111111100000000",
				"0000000000000000111111100000000",
				"0000000000000000111111100000000",
				"0000000000000000111111100000000",
				"0000000011110000111111100000000",
				"0000000011110000011111100000000",
				"0000000011111000111111100000000",
				"0000000011110000111111000000000",
				"0000000011110000111111000000000",
				"0000000001110000111110000000000",
				"0000000001111001111100000000000",
				"0000000000111111111000000000000",
				"0000000000001111100000000000000",
				"0000000000000000000000000000000"
					);

constant SIX: char:= (
				"0000000000000000000000000000000",
				"0000000000000000111110000000000",
				"0000000000000111111110000000000",
				"0000000000001111111000000000000",
				"0000000000011111000000000000000",
				"0000000000111110000000000000000",
				"0000000001111100000000000000000",
				"0000000001111100000000000000000",
				"0000000011111100000000000000000",
				"0000000011111101111000000000000",
				"0000000011111111111110000000000",
				"0000000011111111111111000000000",
				"0000000111111100111111000000000",
				"0000000111111100011111100000000",
				"0000000111111100011111100000000",
				"0000000111111100011111100000000",
				"0000000111111100011111100000000",
				"0000000111111100011111100000000",
				"0000000111111100011111100000000",
				"0000000111111100011111100000000",
				"0000000111111100011111100000000",
				"0000000111111100011111100000000",
				"0000000011111100011111100000000",
				"0000000011111100011111100000000",
				"0000000011111100011111000000000",
				"0000000011111100011111000000000",
				"0000000001111100011110000000000",
				"0000000000111100111110000000000",
				"0000000000111111111100000000000",
				"0000000000001111110000000000000",
				"0000000000000000000000000000000"
					);
					
constant SEVEN: char:= (
				"0000000000000000000000000000000",
				"0000000011111111111111110000000",
				"0000000011111111111111100000000",
				"0000000011111111111111100000000",
				"0000000011111111111111100000000",
				"0000000011111111111111000000000",
				"0000000011100000000111000000000",
				"0000000011000000000110000000000",
				"0000000010000000001110000000000",
				"0000000000000000001110000000000",
				"0000000000000000011100000000000",
				"0000000000000000111100000000000",
				"0000000000000000111100000000000",
				"0000000000000001111100000000000",
				"0000000000000001111000000000000",
				"0000000000000001111000000000000",
				"0000000000000011111000000000000",
				"0000000000000011111000000000000",
				"0000000000000011111000000000000",
				"0000000000000111111000000000000",
				"0000000000000111111000000000000",
				"0000000000000111111000000000000",
				"0000000000000111111000000000000",
				"0000000000001111111000000000000",
				"0000000000001111111000000000000",
				"0000000000001111111000000000000",
				"0000000000001111111000000000000",
				"0000000000011111111100000000000",
				"0000000000011111111100000000000",
				"0000000000000000000000000000000",
				"0000000000000000000000000000000"
					);

constant EIGHT: char:= (
				"0000000000000000000000000000000",
				"0000000000000111111000000000000",
				"0000000000011111111110000000000",
				"0000000000111110001111000000000",
				"0000000001111100000111000000000",
				"0000000001111000000111100000000",
				"0000000011111000000111100000000",
				"0000000011111000000111100000000",
				"0000000011111100000111100000000",
				"0000000011111110000111100000000",
				"0000000011111111000111000000000",
				"0000000001111111101111000000000",
				"0000000001111111111110000000000",
				"0000000000111111111100000000000",
				"0000000000011111111110000000000",
				"0000000000011111111111000000000",
				"0000000000111111111111000000000",
				"0000000001111011111111100000000",
				"0000000001110001111111100000000",
				"0000000011110000011111110000000",
				"0000000011110000001111110000000",
				"0000000011110000001111110000000",
				"0000000011110000000111110000000",
				"0000000011110000000111100000000",
				"0000000011110000000111100000000",
				"0000000011110000000111100000000",
				"0000000001111000001111000000000",
				"0000000001111100011111000000000",
				"0000000000111111111100000000000",
				"0000000000001111111000000000000",
				"0000000000000000000000000000000"
					);

constant NINE: char:= (
				"0000000000000000000000000000000",
				"0000000000001111100000000000000",
				"0000000000111111111000000000000",
				"0000000001111100111100000000000",
				"0000000001111000111110000000000",
				"0000000011111000111110000000000",
				"0000000011111000111111000000000",
				"0000000111111000111111000000000",
				"0000000111111000111111000000000",
				"0000000111111000111111000000000",
				"0000000111111000111111000000000",
				"0000000111111000111111100000000",
				"0000000111111000111111100000000",
				"0000000111111000111111100000000",
				"0000000111111000111111100000000",
				"0000000111111000111111100000000",
				"0000000111111000111111100000000",
				"0000000111111000111111100000000",
				"0000000011111000111111000000000",
				"0000000011111111111111000000000",
				"0000000001111111111111000000000",
				"0000000000111110111111000000000",
				"0000000000000000111111000000000",
				"0000000000000000111110000000000",
				"0000000000000000111110000000000",
				"0000000000000001111100000000000",
				"0000000000000011111000000000000",
				"0000000000001111110000000000000",
				"0000000001111111100000000000000",
				"0000000001111110000000000000000",
				"0000000000000000000000000000000"
					);

constant V: char:=(
				"0000000000000000000000000000000",
				"0000000000000000000000000000000",
				"0111111111000000000000111111110",
				"0011111111000000000001111111110",
				"0011111111100000000001111111100",
				"0001111111100000000001111111100",
				"0001111111100000000011111111000",
				"0001111111100000000011111111000",
				"0000111111110000000011111111000",
				"0000111111110000000011111110000",
				"0000111111110000000111111110000",
				"0000011111111000000111111110000",
				"0000011111111000000111111100000",
				"0000001111111000001111111100000",
				"0000001111111100001111111000000",
				"0000001111111100001111111000000",
				"0000000111111100011111111000000",
				"0000000111111110011111110000000",
				"0000000111111110011111110000000",
				"0000000011111110111111110000000",
				"0000000011111111111111100000000",
				"0000000001111111111111100000000",
				"0000000001111111111111000000000",
				"0000000001111111111111000000000",
				"0000000000111111111111000000000",
				"0000000000111111111110000000000",
				"0000000000011111111110000000000",
				"0000000000011111111110000000000",
				"0000000000011111111100000000000",
				"0000000000000000000000000000000",
				"0000000000000000000000000000000"
					);
