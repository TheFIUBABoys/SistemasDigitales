-- 67 x 67 px

constant ZERO: char:= (
				"0000000000000000000000000000000000000000000000000000000000000000000",
				"0000000000000000000000000000011110000000000000000000000000000000000",
				"0000000000000000000000000001111111100000000000000000000000000000000",
				"0000000000000000000000000011111111110000000000000000000000000000000",
				"0000000000000000000000000111111111111000000000000000000000000000000",
				"0000000000000000000000001111111111111100000000000000000000000000000",
				"0000000000000000000000011111110011111110000000000000000000000000000",
				"0000000000000000000000011111100001111110000000000000000000000000000",
				"0000000000000000000000111111100001111111000000000000000000000000000",
				"0000000000000000000000111111100001111111000000000000000000000000000",
				"0000000000000000000000111111100001111111000000000000000000000000000",
				"0000000000000000000001111111100001111111100000000000000000000000000",
				"0000000000000000000001111111100001111111100000000000000000000000000",
				"0000000000000000000001111111100001111111100000000000000000000000000",
				"0000000000000000000001111111100001111111110000000000000000000000000",
				"0000000000000000000011111111100001111111110000000000000000000000000",
				"0000000000000000000011111111100001111111110000000000000000000000000",
				"0000000000000000000011111111100001111111110000000000000000000000000",
				"0000000000000000000011111111100001111111111000000000000000000000000",
				"0000000000000000000011111111100001111111111000000000000000000000000",
				"0000000000000000000011111111100001111111111000000000000000000000000",
				"0000000000000000000111111111100001111111111000000000000000000000000",
				"0000000000000000000111111111100001111111111000000000000000000000000",
				"0000000000000000000111111111100001111111111000000000000000000000000",
				"0000000000000000000111111111100001111111111000000000000000000000000",
				"0000000000000000000111111111100001111111111000000000000000000000000",
				"0000000000000000000111111111100001111111111000000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111000000000000000000000000",
				"0000000000000000000111111111100001111111111000000000000000000000000",
				"0000000000000000000111111111100001111111111000000000000000000000000",
				"0000000000000000000111111111100001111111111000000000000000000000000",
				"0000000000000000000111111111100001111111111000000000000000000000000",
				"0000000000000000000111111111100001111111111000000000000000000000000",
				"0000000000000000000111111111100001111111111000000000000000000000000",
				"0000000000000000000011111111100001111111111000000000000000000000000",
				"0000000000000000000011111111100001111111111000000000000000000000000",
				"0000000000000000000011111111100001111111110000000000000000000000000",
				"0000000000000000000011111111100001111111110000000000000000000000000",
				"0000000000000000000011111111100001111111110000000000000000000000000",
				"0000000000000000000001111111100001111111110000000000000000000000000",
				"0000000000000000000001111111100001111111100000000000000000000000000",
				"0000000000000000000001111111100001111111100000000000000000000000000",
				"0000000000000000000001111111100001111111100000000000000000000000000",
				"0000000000000000000000111111100001111111100000000000000000000000000",
				"0000000000000000000000111111100001111111000000000000000000000000000",
				"0000000000000000000000011111100001111111000000000000000000000000000",
				"0000000000000000000000011111100001111110000000000000000000000000000",
				"0000000000000000000000001111110001111110000000000000000000000000000",
				"0000000000000000000000001111111111111100000000000000000000000000000",
				"0000000000000000000000000111111111111000000000000000000000000000000",
				"0000000000000000000000000011111111110000000000000000000000000000000",
				"0000000000000000000000000001111111100000000000000000000000000000000",
				"0000000000000000000000000000111111000000000000000000000000000000000",
				"0000000000000000000000000000000000000000000000000000000000000000000"
					);
					
constant ONE: char:= (
				"000000000000000000000000000000000000000000000000000000000000000000000",
				"000000000000000000000000000000000000011100000000000000000000000000000",
				"000000000000000000000000000000000000111100000000000000000000000000000",
				"000000000000000000000000000000000001111100000000000000000000000000000",
				"000000000000000000000000000000000001111100000000000000000000000000000",
				"000000000000000000000000000000000011111100000000000000000000000000000",
				"000000000000000000000000000000000011111100000000000000000000000000000",
				"000000000000000000000000000000000111111100000000000000000000000000000",
				"000000000000000000000000000000000111111100000000000000000000000000000",
				"000000000000000000000000000000001111111100000000000000000000000000000",
				"000000000000000000000000000000011111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000001111111111100000000000000000000000000000",
				"000000000000000000000000000011111111111100000000000000000000000000000",
				"000000000000000000000000000111111111111100000000000000000000000000000",
				"000000000000000000000000001111111111111100000000000000000000000000000",
				"000000000000000000000000011111111111111100000000000000000000000000000",
				"000000000000000000000000011111111111111100000000000000000000000000000",
				"000000000000000000000000011111111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000000111111111100000000000000000000000000000",
				"000000000000000000000000000011111111111110000000000000000000000000000",
				"000000000000000000000000000011111111111111000000000000000000000000000",
				"000000000000000000000000000011111111111111000000000000000000000000000",
				"000000000000000000000000000011111111111111000000000000000000000000000",
				"000000000000000000000000000011111111111111000000000000000000000000000",
				"000000000000000000000000000011111111111111000000000000000000000000000",
				"000000000000000000000000000000000000000000000000000000000000000000000"
					);

constant TWO: char:= (
				"0000000000000000000000000000000000000000000000000000000000000000000",
				"0000000000000000000000000000001111100000000000000000000000000000000",
				"0000000000000000000000000001111111111100000000000000000000000000000",
				"0000000000000000000000000011111111111110000000000000000000000000000",
				"0000000000000000000000000111111111111111000000000000000000000000000",
				"0000000000000000000000001111111111111111100000000000000000000000000",
				"0000000000000000000000011111110001111111110000000000000000000000000",
				"0000000000000000000000011111100000111111110000000000000000000000000",
				"0000000000000000000000111111100000111111111000000000000000000000000",
				"0000000000000000000000111111000000111111111000000000000000000000000",
				"0000000000000000000000111111000000011111111100000000000000000000000",
				"0000000000000000000001111111000000011111111100000000000000000000000",
				"0000000000000000000001111111100000011111111100000000000000000000000",
				"0000000000000000000001111111100000011111111110000000000000000000000",
				"0000000000000000000001111111100000011111111110000000000000000000000",
				"0000000000000000000001111111100000011111111110000000000000000000000",
				"0000000000000000000001111111100000011111111110000000000000000000000",
				"0000000000000000000001111111100000011111111110000000000000000000000",
				"0000000000000000000001111111000000011111111110000000000000000000000",
				"0000000000000000000001111111000000011111111110000000000000000000000",
				"0000000000000000000000111111000000011111111110000000000000000000000",
				"0000000000000000000000111110000000011111111110000000000000000000000",
				"0000000000000000000000011110000000011111111110000000000000000000000",
				"0000000000000000000000000000000000011111111110000000000000000000000",
				"0000000000000000000000000000000000011111111110000000000000000000000",
				"0000000000000000000000000000000000111111111100000000000000000000000",
				"0000000000000000000000000000000000111111111100000000000000000000000",
				"0000000000000000000000000000000000111111111100000000000000000000000",
				"0000000000000000000000000000000000111111111100000000000000000000000",
				"0000000000000000000000000000000000111111111000000000000000000000000",
				"0000000000000000000000000000000001111111111000000000000000000000000",
				"0000000000000000000000000000000001111111110000000000000000000000000",
				"0000000000000000000000000000000001111111110000000000000000000000000",
				"0000000000000000000000000000000011111111100000000000000000000000000",
				"0000000000000000000000000000000011111111100000000000000000000000000",
				"0000000000000000000000000000000011111111000000000000000000000000000",
				"0000000000000000000000000000000111111110000000000000000000000000000",
				"0000000000000000000000000000000111111100000000000000000000000000000",
				"0000000000000000000000000000001111111100000000000000000000000000000",
				"0000000000000000000000000000001111111000000000000000000000000000000",
				"0000000000000000000000000000011111110000000000000000000000000000000",
				"0000000000000000000000000000011111100000000000000000000000000000000",
				"0000000000000000000000000000111111000000000000000000000000000000000",
				"0000000000000000000000000001111110000000000000000000000000000000000",
				"0000000000000000000000000001111110000000000000000000000000000000000",
				"0000000000000000000000000011111100000000000000000000000000000000000",
				"0000000000000000000000000011111000000000000000000000000000000000000",
				"0000000000000000000000000111110000000000001110000000000000000000000",
				"0000000000000000000000000111100000000000001110000000000000000000000",
				"0000000000000000000000001111100000000000001110000000000000000000000",
				"0000000000000000000000011111000000000000001110000000000000000000000",
				"0000000000000000000000011110000000000000001110000000000000000000000",
				"0000000000000000000000111100000000000000011110000000000000000000000",
				"0000000000000000000001111100000000000000011110000000000000000000000",
				"0000000000000000000001111111111111111111111110000000000000000000000",
				"0000000000000000000001111111111111111111111110000000000000000000000",
				"0000000000000000000001111111111111111111111110000000000000000000000",
				"0000000000000000000001111111111111111111111100000000000000000000000",
				"0000000000000000000001111111111111111111111100000000000000000000000",
				"0000000000000000000001111111111111111111111100000000000000000000000",
				"0000000000000000000001111111111111111111111100000000000000000000000",
				"0000000000000000000001111111111111111111111100000000000000000000000",
				"0000000000000000000001111111111111111111111100000000000000000000000",
				"0000000000000000000001111111111111111111111100000000000000000000000",
				"0000000000000000000001111111111111111111111000000000000000000000000",
				"0000000000000000000001111111111111111111111000000000000000000000000",
				"0000000000000000000000000000000000000000000000000000000000000000000"
					);

constant THREE: char:= (
				"0000000000000000000000000000000000000000000000000000000000000000000",
				"0000000000000000000000000000111111111000000000000000000000000000000",
				"0000000000000000000000000001111111111110000000000000000000000000000",
				"0000000000000000000000000011111111111111000000000000000000000000000",
				"0000000000000000000000000111111111111111100000000000000000000000000",
				"0000000000000000000000001111111111111111100000000000000000000000000",
				"0000000000000000000000001111100001111111110000000000000000000000000",
				"0000000000000000000000011111100001111111110000000000000000000000000",
				"0000000000000000000000011111000000111111111000000000000000000000000",
				"0000000000000000000000111111000000111111111000000000000000000000000",
				"0000000000000000000000111111000000111111111000000000000000000000000",
				"0000000000000000000000111111100000111111111100000000000000000000000",
				"0000000000000000000000111111100000111111111100000000000000000000000",
				"0000000000000000000000111111100000111111111100000000000000000000000",
				"0000000000000000000000111111100000111111111100000000000000000000000",
				"0000000000000000000000111111100000111111111100000000000000000000000",
				"0000000000000000000000111111100000111111111100000000000000000000000",
				"0000000000000000000000111111100000111111111100000000000000000000000",
				"0000000000000000000000011111100000111111111100000000000000000000000",
				"0000000000000000000000011111000000111111111100000000000000000000000",
				"0000000000000000000000001111000000111111111100000000000000000000000",
				"0000000000000000000000000000000000111111111100000000000000000000000",
				"0000000000000000000000000000000000111111111000000000000000000000000",
				"0000000000000000000000000000000000111111111000000000000000000000000",
				"0000000000000000000000000000000000111111110000000000000000000000000",
				"0000000000000000000000000000000000111111110000000000000000000000000",
				"0000000000000000000000000000000001111111100000000000000000000000000",
				"0000000000000000000000000000000011111111100000000000000000000000000",
				"0000000000000000000000000000001111111111000000000000000000000000000",
				"0000000000000000000000000011111111111100000000000000000000000000000",
				"0000000000000000000000000011111111110000000000000000000000000000000",
				"0000000000000000000000000011111111110000000000000000000000000000000",
				"0000000000000000000000000011111111111100000000000000000000000000000",
				"0000000000000000000000000011111111111111000000000000000000000000000",
				"0000000000000000000000000000000011111111100000000000000000000000000",
				"0000000000000000000000000000000001111111110000000000000000000000000",
				"0000000000000000000000000000000000111111110000000000000000000000000",
				"0000000000000000000000000000000000111111111000000000000000000000000",
				"0000000000000000000000000000000000111111111100000000000000000000000",
				"0000000000000000000000000000000000111111111100000000000000000000000",
				"0000000000000000000000000000000000111111111100000000000000000000000",
				"0000000000000000000000000000000000011111111110000000000000000000000",
				"0000000000000000000000000000000000011111111110000000000000000000000",
				"0000000000000000000000000000000000011111111110000000000000000000000",
				"0000000000000000000000000000000000011111111110000000000000000000000",
				"0000000000000000000000001100000000011111111110000000000000000000000",
				"0000000000000000000000011111000000011111111110000000000000000000000",
				"0000000000000000000000111111000000011111111110000000000000000000000",
				"0000000000000000000000111111000000011111111110000000000000000000000",
				"0000000000000000000000111111100000011111111110000000000000000000000",
				"0000000000000000000001111111100000011111111110000000000000000000000",
				"0000000000000000000001111111100000011111111110000000000000000000000",
				"0000000000000000000001111111100000011111111110000000000000000000000",
				"0000000000000000000001111111100000011111111110000000000000000000000",
				"0000000000000000000000111111100000011111111100000000000000000000000",
				"0000000000000000000000111111000000011111111100000000000000000000000",
				"0000000000000000000000111111000000011111111100000000000000000000000",
				"0000000000000000000000111111000000111111111000000000000000000000000",
				"0000000000000000000000011111000000111111111000000000000000000000000",
				"0000000000000000000000011111100000111111110000000000000000000000000",
				"0000000000000000000000011111100001111111110000000000000000000000000",
				"0000000000000000000000001111111111111111100000000000000000000000000",
				"0000000000000000000000000111111111111111000000000000000000000000000",
				"0000000000000000000000000011111111111110000000000000000000000000000",
				"0000000000000000000000000001111111111100000000000000000000000000000",
				"0000000000000000000000000000111111110000000000000000000000000000000",
				"0000000000000000000000000000000000000000000000000000000000000000000"
					);

constant FOUR: char:= (
				"0000000000000000000000000000000000000000000000000000000000000000000",
				"0000000000000000000000000000000000001111000000000000000000000000000",
				"0000000000000000000000000000000000011111000000000000000000000000000",
				"0000000000000000000000000000000000011111000000000000000000000000000",
				"0000000000000000000000000000000000011111000000000000000000000000000",
				"0000000000000000000000000000000000111111000000000000000000000000000",
				"0000000000000000000000000000000000111111000000000000000000000000000",
				"0000000000000000000000000000000001111111000000000000000000000000000",
				"0000000000000000000000000000000001111111000000000000000000000000000",
				"0000000000000000000000000000000011111111000000000000000000000000000",
				"0000000000000000000000000000000011111111000000000000000000000000000",
				"0000000000000000000000000000000011111111000000000000000000000000000",
				"0000000000000000000000000000000111111111000000000000000000000000000",
				"0000000000000000000000000000000111111111000000000000000000000000000",
				"0000000000000000000000000000001111111111000000000000000000000000000",
				"0000000000000000000000000000001111111111000000000000000000000000000",
				"0000000000000000000000000000011111111111000000000000000000000000000",
				"0000000000000000000000000000011111111111000000000000000000000000000",
				"0000000000000000000000000000111111111111000000000000000000000000000",
				"0000000000000000000000000000111111111111000000000000000000000000000",
				"0000000000000000000000000000111111111111000000000000000000000000000",
				"0000000000000000000000000001111111111111000000000000000000000000000",
				"0000000000000000000000000001111111111111000000000000000000000000000",
				"0000000000000000000000000011110111111111000000000000000000000000000",
				"0000000000000000000000000011110111111111000000000000000000000000000",
				"0000000000000000000000000111100111111111000000000000000000000000000",
				"0000000000000000000000000111100111111111000000000000000000000000000",
				"0000000000000000000000000111000111111111000000000000000000000000000",
				"0000000000000000000000001111000111111111000000000000000000000000000",
				"0000000000000000000000001111000111111111000000000000000000000000000",
				"0000000000000000000000011110000111111111000000000000000000000000000",
				"0000000000000000000000011110000111111111000000000000000000000000000",
				"0000000000000000000000111100000111111111000000000000000000000000000",
				"0000000000000000000000111100000111111111000000000000000000000000000",
				"0000000000000000000000111000000111111111000000000000000000000000000",
				"0000000000000000000001111000000111111111000000000000000000000000000",
				"0000000000000000000001111000000111111111000000000000000000000000000",
				"0000000000000000000011110000000111111111000000000000000000000000000",
				"0000000000000000000011110000000111111111000000000000000000000000000",
				"0000000000000000000111100000000111111111000000000000000000000000000",
				"0000000000000000000111100000000111111111000000000000000000000000000",
				"0000000000000000000111000000000111111111000000000000000000000000000",
				"0000000000000000000111000000000111111111000000000000000000000000000",
				"0000000000000000000111111111111111111111111100000000000000000000000",
				"0000000000000000000111111111111111111111111100000000000000000000000",
				"0000000000000000000111111111111111111111111100000000000000000000000",
				"0000000000000000000111111111111111111111111100000000000000000000000",
				"0000000000000000000111111111111111111111111100000000000000000000000",
				"0000000000000000000111111111111111111111111100000000000000000000000",
				"0000000000000000000000000000000111111111000000000000000000000000000",
				"0000000000000000000000000000000111111111000000000000000000000000000",
				"0000000000000000000000000000000111111111000000000000000000000000000",
				"0000000000000000000000000000000111111111000000000000000000000000000",
				"0000000000000000000000000000000111111111000000000000000000000000000",
				"0000000000000000000000000000000111111111000000000000000000000000000",
				"0000000000000000000000000000000111111111000000000000000000000000000",
				"0000000000000000000000000000000111111111000000000000000000000000000",
				"0000000000000000000000000000000111111111000000000000000000000000000",
				"0000000000000000000000000000000111111111000000000000000000000000000",
				"0000000000000000000000000000001111111111100000000000000000000000000",
				"0000000000000000000000000000001111111111110000000000000000000000000",
				"0000000000000000000000000000011111111111110000000000000000000000000",
				"0000000000000000000000000000011111111111110000000000000000000000000",
				"0000000000000000000000000000011111111111110000000000000000000000000",
				"0000000000000000000000000000011111111111110000000000000000000000000",
				"0000000000000000000000000000011111111111110000000000000000000000000",
				"0000000000000000000000000000000000000000000000000000000000000000000"
					);

constant FIVE: char:= (
				"0000000000000000000000000000000000000000000000000000000000000000000",
				"0000000000000000000000000000000000000011100000000000000000000000000",
				"0000000000000000000000001111111111111111100000000000000000000000000",
				"0000000000000000000000011111111111111111100000000000000000000000000",
				"0000000000000000000000011111111111111111100000000000000000000000000",
				"0000000000000000000000011111111111111111100000000000000000000000000",
				"0000000000000000000000011111111111111111100000000000000000000000000",
				"0000000000000000000000011111111111111111100000000000000000000000000",
				"0000000000000000000000011111111111111111100000000000000000000000000",
				"0000000000000000000000011111111111111111100000000000000000000000000",
				"0000000000000000000000011111111111111111000000000000000000000000000",
				"0000000000000000000000011111111111111111000000000000000000000000000",
				"0000000000000000000000011111111111111111000000000000000000000000000",
				"0000000000000000000000011111111111111111000000000000000000000000000",
				"0000000000000000000000011100000000000000000000000000000000000000000",
				"0000000000000000000000011100000000000000000000000000000000000000000",
				"0000000000000000000000011100000000000000000000000000000000000000000",
				"0000000000000000000000011100000000000000000000000000000000000000000",
				"0000000000000000000000011100000000000000000000000000000000000000000",
				"0000000000000000000000011100000000000000000000000000000000000000000",
				"0000000000000000000000011100000000000000000000000000000000000000000",
				"0000000000000000000000011100000000000000000000000000000000000000000",
				"0000000000000000000000011100000000000000000000000000000000000000000",
				"0000000000000000000000011100000000000000000000000000000000000000000",
				"0000000000000000000000011100111111110000000000000000000000000000000",
				"0000000000000000000000111101111111111000000000000000000000000000000",
				"0000000000000000000000111111111111111110000000000000000000000000000",
				"0000000000000000000000111111111111111110000000000000000000000000000",
				"0000000000000000000000111111111111111111000000000000000000000000000",
				"0000000000000000000000111111000111111111100000000000000000000000000",
				"0000000000000000000000111110000011111111100000000000000000000000000",
				"0000000000000000000000111110000001111111110000000000000000000000000",
				"0000000000000000000000111100000001111111110000000000000000000000000",
				"0000000000000000000000111100000001111111111000000000000000000000000",
				"0000000000000000000000111100000001111111111000000000000000000000000",
				"0000000000000000000000111000000001111111111000000000000000000000000",
				"0000000000000000000000000000000000111111111000000000000000000000000",
				"0000000000000000000000000000000000111111111100000000000000000000000",
				"0000000000000000000000000000000000111111111100000000000000000000000",
				"0000000000000000000000000000000000111111111100000000000000000000000",
				"0000000000000000000000000000000000111111111100000000000000000000000",
				"0000000000000000000000000000000000111111111100000000000000000000000",
				"0000000000000000000000000000000000111111111100000000000000000000000",
				"0000000000000000000000000000000000111111111100000000000000000000000",
				"0000000000000000000000000000000000111111111100000000000000000000000",
				"0000000000000000000000000000000000111111111100000000000000000000000",
				"0000000000000000000000111100000000111111111100000000000000000000000",
				"0000000000000000000000111110000000111111111100000000000000000000000",
				"0000000000000000000001111110000000111111111100000000000000000000000",
				"0000000000000000000001111110000000111111111100000000000000000000000",
				"0000000000000000000011111110000000111111111100000000000000000000000",
				"0000000000000000000011111111000000111111111100000000000000000000000",
				"0000000000000000000011111111000000111111111000000000000000000000000",
				"0000000000000000000011111110000000111111111000000000000000000000000",
				"0000000000000000000011111110000000111111111000000000000000000000000",
				"0000000000000000000011111110000000111111111000000000000000000000000",
				"0000000000000000000001111110000000111111110000000000000000000000000",
				"0000000000000000000001111110000000111111110000000000000000000000000",
				"0000000000000000000001111110000001111111100000000000000000000000000",
				"0000000000000000000000111110000001111111100000000000000000000000000",
				"0000000000000000000000111111000011111111000000000000000000000000000",
				"0000000000000000000000011111100111111110000000000000000000000000000",
				"0000000000000000000000011111111111111110000000000000000000000000000",
				"0000000000000000000000001111111111111100000000000000000000000000000",
				"0000000000000000000000000111111111110000000000000000000000000000000",
				"0000000000000000000000000011111111100000000000000000000000000000000",
				"0000000000000000000000000000000000000000000000000000000000000000000"
					);

constant SIX: char:= (
				"0000000000000000000000000000000000000000000000000000000000000000000",
				"0000000000000000000000000000000000001111100000000000000000000000000",
				"0000000000000000000000000000000001111111100000000000000000000000000",
				"0000000000000000000000000000000111111111100000000000000000000000000",
				"0000000000000000000000000000001111111111100000000000000000000000000",
				"0000000000000000000000000000111111111111100000000000000000000000000",
				"0000000000000000000000000001111111111110000000000000000000000000000",
				"0000000000000000000000000011111111110000000000000000000000000000000",
				"0000000000000000000000000011111111000000000000000000000000000000000",
				"0000000000000000000000000111111110000000000000000000000000000000000",
				"0000000000000000000000001111111100000000000000000000000000000000000",
				"0000000000000000000000001111111100000000000000000000000000000000000",
				"0000000000000000000000011111111000000000000000000000000000000000000",
				"0000000000000000000000011111111000000000000000000000000000000000000",
				"0000000000000000000000011111110000000000000000000000000000000000000",
				"0000000000000000000000111111110000000000000000000000000000000000000",
				"0000000000000000000000111111110000000000000000000000000000000000000",
				"0000000000000000000000111111110000000000000000000000000000000000000",
				"0000000000000000000001111111110000000000000000000000000000000000000",
				"0000000000000000000001111111110001111000000000000000000000000000000",
				"0000000000000000000001111111110011111110000000000000000000000000000",
				"0000000000000000000001111111110111111111000000000000000000000000000",
				"0000000000000000000001111111111111111111100000000000000000000000000",
				"0000000000000000000011111111111111111111100000000000000000000000000",
				"0000000000000000000011111111111111111111110000000000000000000000000",
				"0000000000000000000011111111111101111111110000000000000000000000000",
				"0000000000000000000011111111111000111111111000000000000000000000000",
				"0000000000000000000011111111110000111111111000000000000000000000000",
				"0000000000000000000011111111110000111111111000000000000000000000000",
				"0000000000000000000011111111110000111111111000000000000000000000000",
				"0000000000000000000011111111110000111111111100000000000000000000000",
				"0000000000000000000011111111110000111111111100000000000000000000000",
				"0000000000000000000011111111110000111111111100000000000000000000000",
				"0000000000000000000011111111110000111111111100000000000000000000000",
				"0000000000000000000011111111110000111111111100000000000000000000000",
				"0000000000000000000011111111110000111111111100000000000000000000000",
				"0000000000000000000011111111110000111111111100000000000000000000000",
				"0000000000000000000011111111110000111111111110000000000000000000000",
				"0000000000000000000011111111110000111111111110000000000000000000000",
				"0000000000000000000011111111110000111111111110000000000000000000000",
				"0000000000000000000011111111110000111111111110000000000000000000000",
				"0000000000000000000011111111110000111111111110000000000000000000000",
				"0000000000000000000011111111110000111111111110000000000000000000000",
				"0000000000000000000011111111110000111111111110000000000000000000000",
				"0000000000000000000011111111110000111111111110000000000000000000000",
				"0000000000000000000011111111110000111111111100000000000000000000000",
				"0000000000000000000011111111110000111111111100000000000000000000000",
				"0000000000000000000011111111110000111111111100000000000000000000000",
				"0000000000000000000011111111110000111111111100000000000000000000000",
				"0000000000000000000011111111110000111111111100000000000000000000000",
				"0000000000000000000011111111110000111111111100000000000000000000000",
				"0000000000000000000001111111110000111111111100000000000000000000000",
				"0000000000000000000001111111110000111111111000000000000000000000000",
				"0000000000000000000001111111110000111111111000000000000000000000000",
				"0000000000000000000001111111110000111111111000000000000000000000000",
				"0000000000000000000000111111110000111111111000000000000000000000000",
				"0000000000000000000000111111110000111111110000000000000000000000000",
				"0000000000000000000000111111110000111111110000000000000000000000000",
				"0000000000000000000000011111110000111111100000000000000000000000000",
				"0000000000000000000000011111110000111111100000000000000000000000000",
				"0000000000000000000000001111110000111111000000000000000000000000000",
				"0000000000000000000000001111111001111111000000000000000000000000000",
				"0000000000000000000000000111111111111110000000000000000000000000000",
				"0000000000000000000000000011111111111100000000000000000000000000000",
				"0000000000000000000000000001111111111000000000000000000000000000000",
				"0000000000000000000000000000111111110000000000000000000000000000000",
				"0000000000000000000000000000000000000000000000000000000000000000000"
					);
					
constant SEVEN: char:= (
				"0000000000000000000000000000000000000000000000000000000000000000000",
				"0000000000000000000001111111111111111111111100000000000000000000000",
				"0000000000000000000001111111111111111111111100000000000000000000000",
				"0000000000000000000001111111111111111111111100000000000000000000000",
				"0000000000000000000001111111111111111111111100000000000000000000000",
				"0000000000000000000001111111111111111111111100000000000000000000000",
				"0000000000000000000001111111111111111111111100000000000000000000000",
				"0000000000000000000001111111111111111111111000000000000000000000000",
				"0000000000000000000001111111111111111111111000000000000000000000000",
				"0000000000000000000011111111111111111111111000000000000000000000000",
				"0000000000000000000011111111111111111111110000000000000000000000000",
				"0000000000000000000011111111111111111111110000000000000000000000000",
				"0000000000000000000011111111111111111111110000000000000000000000000",
				"0000000000000000000011111000000000000011110000000000000000000000000",
				"0000000000000000000011110000000000000111100000000000000000000000000",
				"0000000000000000000011110000000000000111100000000000000000000000000",
				"0000000000000000000011110000000000000111100000000000000000000000000",
				"0000000000000000000011100000000000001111100000000000000000000000000",
				"0000000000000000000000000000000000001111000000000000000000000000000",
				"0000000000000000000000000000000000011111000000000000000000000000000",
				"0000000000000000000000000000000000011111000000000000000000000000000",
				"0000000000000000000000000000000000011111000000000000000000000000000",
				"0000000000000000000000000000000000111111000000000000000000000000000",
				"0000000000000000000000000000000000111110000000000000000000000000000",
				"0000000000000000000000000000000000111110000000000000000000000000000",
				"0000000000000000000000000000000001111110000000000000000000000000000",
				"0000000000000000000000000000000001111110000000000000000000000000000",
				"0000000000000000000000000000000011111110000000000000000000000000000",
				"0000000000000000000000000000000011111100000000000000000000000000000",
				"0000000000000000000000000000000011111100000000000000000000000000000",
				"0000000000000000000000000000000011111100000000000000000000000000000",
				"0000000000000000000000000000000111111100000000000000000000000000000",
				"0000000000000000000000000000000111111100000000000000000000000000000",
				"0000000000000000000000000000000111111100000000000000000000000000000",
				"0000000000000000000000000000001111111000000000000000000000000000000",
				"0000000000000000000000000000001111111000000000000000000000000000000",
				"0000000000000000000000000000001111111000000000000000000000000000000",
				"0000000000000000000000000000001111111000000000000000000000000000000",
				"0000000000000000000000000000011111111000000000000000000000000000000",
				"0000000000000000000000000000011111111000000000000000000000000000000",
				"0000000000000000000000000000011111111000000000000000000000000000000",
				"0000000000000000000000000000011111111000000000000000000000000000000",
				"0000000000000000000000000000011111111000000000000000000000000000000",
				"0000000000000000000000000000111111111000000000000000000000000000000",
				"0000000000000000000000000000111111111000000000000000000000000000000",
				"0000000000000000000000000000111111111000000000000000000000000000000",
				"0000000000000000000000000000111111111000000000000000000000000000000",
				"0000000000000000000000000000111111111000000000000000000000000000000",
				"0000000000000000000000000000111111111000000000000000000000000000000",
				"0000000000000000000000000001111111111000000000000000000000000000000",
				"0000000000000000000000000001111111111000000000000000000000000000000",
				"0000000000000000000000000001111111111000000000000000000000000000000",
				"0000000000000000000000000001111111111000000000000000000000000000000",
				"0000000000000000000000000001111111111000000000000000000000000000000",
				"0000000000000000000000000001111111111000000000000000000000000000000",
				"0000000000000000000000000001111111111000000000000000000000000000000",
				"0000000000000000000000000001111111111000000000000000000000000000000",
				"0000000000000000000000000001111111111000000000000000000000000000000",
				"0000000000000000000000000001111111111000000000000000000000000000000",
				"0000000000000000000000000011111111111100000000000000000000000000000",
				"0000000000000000000000000111111111111100000000000000000000000000000",
				"0000000000000000000000000111111111111110000000000000000000000000000",
				"0000000000000000000000000111111111111110000000000000000000000000000",
				"0000000000000000000000000111111111111110000000000000000000000000000",
				"0000000000000000000000000011111111111100000000000000000000000000000",
				"0000000000000000000000000000000000000000000000000000000000000000000",
				"0000000000000000000000000000000000000000000000000000000000000000000"
					);

constant EIGHT: char:= (
				"0000000000000000000000000000000000000000000000000000000000000000000",
				"0000000000000000000000000000001111000000000000000000000000000000000",
				"0000000000000000000000000001111111111000000000000000000000000000000",
				"0000000000000000000000000011111111111110000000000000000000000000000",
				"0000000000000000000000000111111111111111000000000000000000000000000",
				"0000000000000000000000001111111111111111000000000000000000000000000",
				"0000000000000000000000011111111000111111100000000000000000000000000",
				"0000000000000000000000011111110000001111110000000000000000000000000",
				"0000000000000000000000111111100000001111110000000000000000000000000",
				"0000000000000000000000111111100000000111110000000000000000000000000",
				"0000000000000000000001111111000000000111111000000000000000000000000",
				"0000000000000000000001111111000000000111111000000000000000000000000",
				"0000000000000000000001111111000000000011111000000000000000000000000",
				"0000000000000000000001111111000000000011111000000000000000000000000",
				"0000000000000000000001111111000000000011111000000000000000000000000",
				"0000000000000000000001111111000000000011111000000000000000000000000",
				"0000000000000000000011111111000000000011111000000000000000000000000",
				"0000000000000000000011111111100000000011111000000000000000000000000",
				"0000000000000000000011111111100000000011111000000000000000000000000",
				"0000000000000000000001111111110000000011111000000000000000000000000",
				"0000000000000000000001111111110000000111111000000000000000000000000",
				"0000000000000000000001111111111000000111111000000000000000000000000",
				"0000000000000000000001111111111100000111110000000000000000000000000",
				"0000000000000000000001111111111110000111110000000000000000000000000",
				"0000000000000000000001111111111111001111100000000000000000000000000",
				"0000000000000000000000111111111111111111100000000000000000000000000",
				"0000000000000000000000111111111111111111000000000000000000000000000",
				"0000000000000000000000111111111111111110000000000000000000000000000",
				"0000000000000000000000011111111111111100000000000000000000000000000",
				"0000000000000000000000011111111111111110000000000000000000000000000",
				"0000000000000000000000001111111111111110000000000000000000000000000",
				"0000000000000000000000001111111111111111000000000000000000000000000",
				"0000000000000000000000000111111111111111100000000000000000000000000",
				"0000000000000000000000000011111111111111100000000000000000000000000",
				"0000000000000000000000000111111111111111110000000000000000000000000",
				"0000000000000000000000001111111111111111110000000000000000000000000",
				"0000000000000000000000011111111111111111111000000000000000000000000",
				"0000000000000000000000111110011111111111111000000000000000000000000",
				"0000000000000000000000111110001111111111111000000000000000000000000",
				"0000000000000000000001111110000111111111111100000000000000000000000",
				"0000000000000000000001111100000011111111111100000000000000000000000",
				"0000000000000000000001111100000001111111111100000000000000000000000",
				"0000000000000000000011111100000001111111111100000000000000000000000",
				"0000000000000000000011111100000000111111111100000000000000000000000",
				"0000000000000000000011111100000000011111111100000000000000000000000",
				"0000000000000000000011111100000000011111111100000000000000000000000",
				"0000000000000000000011111100000000001111111100000000000000000000000",
				"0000000000000000000011111100000000000111111100000000000000000000000",
				"0000000000000000000011111100000000000111111100000000000000000000000",
				"0000000000000000000011111100000000000111111100000000000000000000000",
				"0000000000000000000011111100000000000111111100000000000000000000000",
				"0000000000000000000011111100000000000111111100000000000000000000000",
				"0000000000000000000011111100000000000111111100000000000000000000000",
				"0000000000000000000011111100000000000111111100000000000000000000000",
				"0000000000000000000011111100000000000111111000000000000000000000000",
				"0000000000000000000011111100000000000111111000000000000000000000000",
				"0000000000000000000001111110000000000111111000000000000000000000000",
				"0000000000000000000001111110000000001111110000000000000000000000000",
				"0000000000000000000001111110000000001111110000000000000000000000000",
				"0000000000000000000000111111000000011111100000000000000000000000000",
				"0000000000000000000000111111100000111111100000000000000000000000000",
				"0000000000000000000000011111111111111111000000000000000000000000000",
				"0000000000000000000000001111111111111110000000000000000000000000000",
				"0000000000000000000000000111111111111100000000000000000000000000000",
				"0000000000000000000000000011111111111000000000000000000000000000000",
				"0000000000000000000000000001111111110000000000000000000000000000000",
				"0000000000000000000000000000000000000000000000000000000000000000000"
					);

constant NINE: char:= (
				"0000000000000000000000000000000000000000000000000000000000000000000",
				"0000000000000000000000000000001110000000000000000000000000000000000",
				"0000000000000000000000000001111111100000000000000000000000000000000",
				"0000000000000000000000000011111111111000000000000000000000000000000",
				"0000000000000000000000000111111111111100000000000000000000000000000",
				"0000000000000000000000001111111111111110000000000000000000000000000",
				"0000000000000000000000011111110011111110000000000000000000000000000",
				"0000000000000000000000011111100001111111000000000000000000000000000",
				"0000000000000000000000111111100001111111000000000000000000000000000",
				"0000000000000000000000111111100001111111100000000000000000000000000",
				"0000000000000000000001111111100001111111100000000000000000000000000",
				"0000000000000000000001111111100001111111110000000000000000000000000",
				"0000000000000000000001111111100001111111110000000000000000000000000",
				"0000000000000000000011111111100001111111110000000000000000000000000",
				"0000000000000000000011111111100001111111110000000000000000000000000",
				"0000000000000000000011111111100001111111111000000000000000000000000",
				"0000000000000000000011111111100001111111111000000000000000000000000",
				"0000000000000000000111111111100001111111111000000000000000000000000",
				"0000000000000000000111111111100001111111111000000000000000000000000",
				"0000000000000000000111111111100001111111111000000000000000000000000",
				"0000000000000000000111111111100001111111111000000000000000000000000",
				"0000000000000000000111111111100001111111111000000000000000000000000",
				"0000000000000000000111111111100001111111111000000000000000000000000",
				"0000000000000000000111111111100001111111111000000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000111111111100001111111111100000000000000000000000",
				"0000000000000000000011111111100001111111111100000000000000000000000",
				"0000000000000000000011111111100001111111111100000000000000000000000",
				"0000000000000000000011111111100001111111111000000000000000000000000",
				"0000000000000000000011111111100001111111111000000000000000000000000",
				"0000000000000000000001111111110011111111111000000000000000000000000",
				"0000000000000000000001111111111111111111111000000000000000000000000",
				"0000000000000000000000111111111111111111111000000000000000000000000",
				"0000000000000000000000111111111111111111111000000000000000000000000",
				"0000000000000000000000011111111101111111111000000000000000000000000",
				"0000000000000000000000001111111101111111111000000000000000000000000",
				"0000000000000000000000000111111001111111110000000000000000000000000",
				"0000000000000000000000000001100001111111110000000000000000000000000",
				"0000000000000000000000000000000001111111110000000000000000000000000",
				"0000000000000000000000000000000001111111110000000000000000000000000",
				"0000000000000000000000000000000001111111100000000000000000000000000",
				"0000000000000000000000000000000001111111100000000000000000000000000",
				"0000000000000000000000000000000001111111100000000000000000000000000",
				"0000000000000000000000000000000011111111000000000000000000000000000",
				"0000000000000000000000000000000011111111000000000000000000000000000",
				"0000000000000000000000000000000111111110000000000000000000000000000",
				"0000000000000000000000000000000111111110000000000000000000000000000",
				"0000000000000000000000000000001111111100000000000000000000000000000",
				"0000000000000000000000000000011111111000000000000000000000000000000",
				"0000000000000000000000000011111111111000000000000000000000000000000",
				"0000000000000000000000111111111111110000000000000000000000000000000",
				"0000000000000000000000111111111111100000000000000000000000000000000",
				"0000000000000000000000111111111110000000000000000000000000000000000",
				"0000000000000000000000111111111100000000000000000000000000000000000",
				"0000000000000000000000111111110000000000000000000000000000000000000",
				"0000000000000000000000000000000000000000000000000000000000000000000"
					);
