library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all; 

entity bloqueProcesamientoYControl is
     port(
          entradaFlipFlop: in std_logic;
          salidaVGA: in std_logic_vector(14 downto 0);	-- salida VGA (TODO: ver mapeo de pines)
     );
end;


architecture b_arq of bloqueProcesamientoYControl is
begin
    
	
	
end architecture;
